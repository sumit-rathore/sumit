///////////////////////////////////////////////////////////////////////////////
//
//   Icron Technology Corporation - Copyright 2012
//
///////////////////////////////////////////////////////////////////////////////
//
//   Title       :  bootloader.v
//   Created     :  2012-05-15
//   Author      :  keithk
//
///////////////////////////////////////////////////////////////////////////////
//
//   Description :
//
//    bootloader verilog code
//
///////////////////////////////////////////////////////////////////////////////
//
//     $Id: slash.hdr,v 1.4 2009/01/20 19:48:46 keithk Exp $
//
///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////

module bootrom
  (
   input               clk,
   input               rst_n,
   input               en,
   input  wire [08:00] addr,
   output reg  [31:00] data
   );

  always@(posedge clk) begin
    if(en) begin
      case (addr)
$i
        default: data <= 32'b0;
      endcase
    end
  end

endmodule
